library ieee;
use ieee.std_logic_1164.all;
library work;
use work.Gates.all;

entity Zero_Check is
	port(A: in std_logic_vector(15 downto 0);
			y : out std_logic);
end entity Zero_Check;

architecture struct of Zero_Check is
	signal s, t: std_logic;
begin
	s <= A(0);
	inst1: for i in 1 to 15 generate
		or1: OR_2 port map(s, A(i), t);
		s <= t;
	end generate;
	inst2: INVERTER port map(t, s);
	y <= s;
end struct;